** Profile: "SCHEMATIC1-LAB_1_analys"  [ E:\Mach_dien_project\LAB1_project\LAB1_project-PSpiceFiles\SCHEMATIC1\LAB_1_analys.sim ] 

** Creating circuit file "LAB_1_analys.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\23.1.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
